module ALUnor (
    input [31:0] a,
    input [31:0] b,
    output [31:0] result
);
	nor(result[0], a[0], b[0]);
	nor(result[1], a[1], b[1]);
	nor(result[2], a[2], b[2]);
	nor(result[3], a[3], b[3]);
	nor(result[4], a[4], b[4]);
	nor(result[5], a[5], b[5]);
	nor(result[6], a[6], b[6]);
	nor(result[7], a[7], b[7]);
	nor(result[8], a[8], b[8]);
	nor(result[9], a[9], b[9]);
	nor(result[10], a[10], b[10]);
	nor(result[11], a[11], b[11]);
	nor(result[12], a[12], b[12]);
	nor(result[13], a[13], b[13]);
	nor(result[14], a[14], b[14]);
	nor(result[15], a[15], b[15]);
	nor(result[16], a[16], b[16]);
	nor(result[17], a[17], b[17]);
	nor(result[18], a[18], b[18]);
	nor(result[19], a[19], b[19]);
	nor(result[20], a[20], b[20]);
	nor(result[21], a[21], b[21]);
	nor(result[22], a[22], b[22]);
	nor(result[23], a[23], b[23]);
	nor(result[24], a[24], b[24]);
	nor(result[25], a[25], b[25]);
	nor(result[26], a[26], b[26]);
	nor(result[27], a[27], b[27]);
	nor(result[28], a[28], b[28]);
	nor(result[29], a[29], b[29]);
	nor(result[30], a[30], b[30]);
	nor(result[31], a[31], b[31]);
	
endmodule