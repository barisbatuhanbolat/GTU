module ALUand (
    input [31:0] a,
    input [31:0] b,
    output [31:0] result
);
	and(result[0], a[0], b[0]);
	and(result[1], a[1], b[1]);
	and(result[2], a[2], b[2]);
	and(result[3], a[3], b[3]);
	and(result[4], a[4], b[4]);
	and(result[5], a[5], b[5]);
	and(result[6], a[6], b[6]);
	and(result[7], a[7], b[7]);
	and(result[8], a[8], b[8]);
	and(result[9], a[9], b[9]);
	and(result[10], a[10], b[10]);
	and(result[11], a[11], b[11]);
	and(result[12], a[12], b[12]);
	and(result[13], a[13], b[13]);
	and(result[14], a[14], b[14]);
	and(result[15], a[15], b[15]);
	and(result[16], a[16], b[16]);
	and(result[17], a[17], b[17]);
	and(result[18], a[18], b[18]);
	and(result[19], a[19], b[19]);
	and(result[20], a[20], b[20]);
	and(result[21], a[21], b[21]);
	and(result[22], a[22], b[22]);
	and(result[23], a[23], b[23]);
	and(result[24], a[24], b[24]);
	and(result[25], a[25], b[25]);
	and(result[26], a[26], b[26]);
	and(result[27], a[27], b[27]);
	and(result[28], a[28], b[28]);
	and(result[29], a[29], b[29]);
	and(result[30], a[30], b[30]);
	and(result[31], a[31], b[31]);
	
endmodule