module alu(input [31:0] A, input [31:0] B, input [2:0] ALUop, output Result);
	
	
	

endmodule