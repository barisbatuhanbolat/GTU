module ALUless-than (
    input [31:0] a,
    input [31:0] b,
	 output less
);

endmodule
	